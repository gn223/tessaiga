module geethanand();
endmodule
